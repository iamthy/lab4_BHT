
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'hdecd60bd;
    ram_cell[       1] = 32'h0;  // 32'h946c667f;
    ram_cell[       2] = 32'h0;  // 32'hd9c9ebf0;
    ram_cell[       3] = 32'h0;  // 32'ha89764ba;
    ram_cell[       4] = 32'h0;  // 32'hf65a5612;
    ram_cell[       5] = 32'h0;  // 32'hc5e04d4f;
    ram_cell[       6] = 32'h0;  // 32'h9387827e;
    ram_cell[       7] = 32'h0;  // 32'hf4a67d02;
    ram_cell[       8] = 32'h0;  // 32'h10027e72;
    ram_cell[       9] = 32'h0;  // 32'h8d4df16a;
    ram_cell[      10] = 32'h0;  // 32'h264cb0b2;
    ram_cell[      11] = 32'h0;  // 32'h5da8f4b3;
    ram_cell[      12] = 32'h0;  // 32'h3248da30;
    ram_cell[      13] = 32'h0;  // 32'h2d56ac1a;
    ram_cell[      14] = 32'h0;  // 32'h0fe48083;
    ram_cell[      15] = 32'h0;  // 32'h4b38919b;
    ram_cell[      16] = 32'h0;  // 32'hfeb7714a;
    ram_cell[      17] = 32'h0;  // 32'h8abc4c80;
    ram_cell[      18] = 32'h0;  // 32'hfa1bc17c;
    ram_cell[      19] = 32'h0;  // 32'hd9deb48c;
    ram_cell[      20] = 32'h0;  // 32'hca301cb6;
    ram_cell[      21] = 32'h0;  // 32'he4bf6e0e;
    ram_cell[      22] = 32'h0;  // 32'hf77f5062;
    ram_cell[      23] = 32'h0;  // 32'h6dede9a5;
    ram_cell[      24] = 32'h0;  // 32'h9fc239d6;
    ram_cell[      25] = 32'h0;  // 32'hccf02be5;
    ram_cell[      26] = 32'h0;  // 32'h3145f6f2;
    ram_cell[      27] = 32'h0;  // 32'h0aa2f28f;
    ram_cell[      28] = 32'h0;  // 32'hb95bde97;
    ram_cell[      29] = 32'h0;  // 32'hfa214318;
    ram_cell[      30] = 32'h0;  // 32'h1aca6014;
    ram_cell[      31] = 32'h0;  // 32'h72fcab08;
    ram_cell[      32] = 32'h0;  // 32'h60c58eda;
    ram_cell[      33] = 32'h0;  // 32'h2c606906;
    ram_cell[      34] = 32'h0;  // 32'hd58734d3;
    ram_cell[      35] = 32'h0;  // 32'h8eb79f26;
    ram_cell[      36] = 32'h0;  // 32'h80628cd7;
    ram_cell[      37] = 32'h0;  // 32'h96986d91;
    ram_cell[      38] = 32'h0;  // 32'h6b291bd7;
    ram_cell[      39] = 32'h0;  // 32'hadf5e9ed;
    ram_cell[      40] = 32'h0;  // 32'hcc4b44b0;
    ram_cell[      41] = 32'h0;  // 32'h647576ed;
    ram_cell[      42] = 32'h0;  // 32'h349a15e2;
    ram_cell[      43] = 32'h0;  // 32'h6fb63e51;
    ram_cell[      44] = 32'h0;  // 32'h17c182ff;
    ram_cell[      45] = 32'h0;  // 32'h49e357fa;
    ram_cell[      46] = 32'h0;  // 32'h628d3124;
    ram_cell[      47] = 32'h0;  // 32'h58a24eee;
    ram_cell[      48] = 32'h0;  // 32'he689d569;
    ram_cell[      49] = 32'h0;  // 32'h1aa6cb9f;
    ram_cell[      50] = 32'h0;  // 32'h0050fd59;
    ram_cell[      51] = 32'h0;  // 32'ha27ab88d;
    ram_cell[      52] = 32'h0;  // 32'hb6840edf;
    ram_cell[      53] = 32'h0;  // 32'h06ea1b06;
    ram_cell[      54] = 32'h0;  // 32'hd5453caa;
    ram_cell[      55] = 32'h0;  // 32'h1d1e2587;
    ram_cell[      56] = 32'h0;  // 32'hbab8daa8;
    ram_cell[      57] = 32'h0;  // 32'h54aef4b3;
    ram_cell[      58] = 32'h0;  // 32'h5f410d36;
    ram_cell[      59] = 32'h0;  // 32'h7536d275;
    ram_cell[      60] = 32'h0;  // 32'h289f67dd;
    ram_cell[      61] = 32'h0;  // 32'h0d7fba6d;
    ram_cell[      62] = 32'h0;  // 32'h39e1b18a;
    ram_cell[      63] = 32'h0;  // 32'h0e15378c;
    ram_cell[      64] = 32'h0;  // 32'h8257f242;
    ram_cell[      65] = 32'h0;  // 32'h82854630;
    ram_cell[      66] = 32'h0;  // 32'h033c01a0;
    ram_cell[      67] = 32'h0;  // 32'h1a6b852e;
    ram_cell[      68] = 32'h0;  // 32'h4576aec5;
    ram_cell[      69] = 32'h0;  // 32'h000e8ce1;
    ram_cell[      70] = 32'h0;  // 32'h140889b7;
    ram_cell[      71] = 32'h0;  // 32'hbc534041;
    ram_cell[      72] = 32'h0;  // 32'h6cd073ad;
    ram_cell[      73] = 32'h0;  // 32'hb752c8f4;
    ram_cell[      74] = 32'h0;  // 32'hecdb66f3;
    ram_cell[      75] = 32'h0;  // 32'h3157b903;
    ram_cell[      76] = 32'h0;  // 32'h3f8409ca;
    ram_cell[      77] = 32'h0;  // 32'h31670c4c;
    ram_cell[      78] = 32'h0;  // 32'hb2d1e99f;
    ram_cell[      79] = 32'h0;  // 32'h9a9e04ed;
    ram_cell[      80] = 32'h0;  // 32'h666fc70d;
    ram_cell[      81] = 32'h0;  // 32'hf09fa497;
    ram_cell[      82] = 32'h0;  // 32'h6e91290d;
    ram_cell[      83] = 32'h0;  // 32'h33858531;
    ram_cell[      84] = 32'h0;  // 32'h68e231ea;
    ram_cell[      85] = 32'h0;  // 32'h2439cab8;
    ram_cell[      86] = 32'h0;  // 32'h5614d8de;
    ram_cell[      87] = 32'h0;  // 32'h7973f0df;
    ram_cell[      88] = 32'h0;  // 32'h25e851be;
    ram_cell[      89] = 32'h0;  // 32'he9c0b37a;
    ram_cell[      90] = 32'h0;  // 32'h9e06f296;
    ram_cell[      91] = 32'h0;  // 32'hcbfbf147;
    ram_cell[      92] = 32'h0;  // 32'h5dc40a68;
    ram_cell[      93] = 32'h0;  // 32'hb4850d6d;
    ram_cell[      94] = 32'h0;  // 32'h1721f7f9;
    ram_cell[      95] = 32'h0;  // 32'h76c587fa;
    ram_cell[      96] = 32'h0;  // 32'h9b487f4c;
    ram_cell[      97] = 32'h0;  // 32'h44e4bb75;
    ram_cell[      98] = 32'h0;  // 32'h482ecdf0;
    ram_cell[      99] = 32'h0;  // 32'h5f521ce7;
    ram_cell[     100] = 32'h0;  // 32'hd7cda65a;
    ram_cell[     101] = 32'h0;  // 32'h27560c4b;
    ram_cell[     102] = 32'h0;  // 32'heb62ff3c;
    ram_cell[     103] = 32'h0;  // 32'h288b2a83;
    ram_cell[     104] = 32'h0;  // 32'h092a0545;
    ram_cell[     105] = 32'h0;  // 32'h09d278ac;
    ram_cell[     106] = 32'h0;  // 32'h9237a640;
    ram_cell[     107] = 32'h0;  // 32'hd11374d9;
    ram_cell[     108] = 32'h0;  // 32'h5d64b879;
    ram_cell[     109] = 32'h0;  // 32'h3a642928;
    ram_cell[     110] = 32'h0;  // 32'hdc97034f;
    ram_cell[     111] = 32'h0;  // 32'ha3e5dfa1;
    ram_cell[     112] = 32'h0;  // 32'hc81d6cdb;
    ram_cell[     113] = 32'h0;  // 32'hb7b7fb54;
    ram_cell[     114] = 32'h0;  // 32'h1c799bc8;
    ram_cell[     115] = 32'h0;  // 32'h33b91b55;
    ram_cell[     116] = 32'h0;  // 32'hb2e820be;
    ram_cell[     117] = 32'h0;  // 32'h759e50a1;
    ram_cell[     118] = 32'h0;  // 32'h3ee7b65c;
    ram_cell[     119] = 32'h0;  // 32'h33088022;
    ram_cell[     120] = 32'h0;  // 32'h07406972;
    ram_cell[     121] = 32'h0;  // 32'h11fe4f96;
    ram_cell[     122] = 32'h0;  // 32'hfbb07877;
    ram_cell[     123] = 32'h0;  // 32'h4176f1d4;
    ram_cell[     124] = 32'h0;  // 32'h55a0060b;
    ram_cell[     125] = 32'h0;  // 32'hf44e263c;
    ram_cell[     126] = 32'h0;  // 32'h572be9a9;
    ram_cell[     127] = 32'h0;  // 32'hdc818dad;
    ram_cell[     128] = 32'h0;  // 32'hfd4bc455;
    ram_cell[     129] = 32'h0;  // 32'hcdb8b56d;
    ram_cell[     130] = 32'h0;  // 32'he2fea65d;
    ram_cell[     131] = 32'h0;  // 32'h486232f0;
    ram_cell[     132] = 32'h0;  // 32'hcc663dc8;
    ram_cell[     133] = 32'h0;  // 32'h301a9ef8;
    ram_cell[     134] = 32'h0;  // 32'h21a4fc48;
    ram_cell[     135] = 32'h0;  // 32'h57155aab;
    ram_cell[     136] = 32'h0;  // 32'h46c2ea65;
    ram_cell[     137] = 32'h0;  // 32'hae273e40;
    ram_cell[     138] = 32'h0;  // 32'h53f84551;
    ram_cell[     139] = 32'h0;  // 32'h137a86b3;
    ram_cell[     140] = 32'h0;  // 32'h86e7f9a1;
    ram_cell[     141] = 32'h0;  // 32'h9cbe7992;
    ram_cell[     142] = 32'h0;  // 32'hfdabdfa4;
    ram_cell[     143] = 32'h0;  // 32'hcd12e1f2;
    ram_cell[     144] = 32'h0;  // 32'hf5752013;
    ram_cell[     145] = 32'h0;  // 32'hdbff0c94;
    ram_cell[     146] = 32'h0;  // 32'h636089a0;
    ram_cell[     147] = 32'h0;  // 32'hb47ae062;
    ram_cell[     148] = 32'h0;  // 32'hc750328f;
    ram_cell[     149] = 32'h0;  // 32'hd32f2c11;
    ram_cell[     150] = 32'h0;  // 32'hfbcf463a;
    ram_cell[     151] = 32'h0;  // 32'h87cb3bdd;
    ram_cell[     152] = 32'h0;  // 32'he5f4388d;
    ram_cell[     153] = 32'h0;  // 32'h895c0b50;
    ram_cell[     154] = 32'h0;  // 32'h51101ab4;
    ram_cell[     155] = 32'h0;  // 32'h32265c78;
    ram_cell[     156] = 32'h0;  // 32'h7a2a353c;
    ram_cell[     157] = 32'h0;  // 32'hed33979c;
    ram_cell[     158] = 32'h0;  // 32'hf8ab4202;
    ram_cell[     159] = 32'h0;  // 32'h355c6809;
    ram_cell[     160] = 32'h0;  // 32'h3cf911b9;
    ram_cell[     161] = 32'h0;  // 32'hb9f699b6;
    ram_cell[     162] = 32'h0;  // 32'h9f886a16;
    ram_cell[     163] = 32'h0;  // 32'h1780bbdd;
    ram_cell[     164] = 32'h0;  // 32'ha671a037;
    ram_cell[     165] = 32'h0;  // 32'h7949dcf7;
    ram_cell[     166] = 32'h0;  // 32'h3107c90d;
    ram_cell[     167] = 32'h0;  // 32'hc2798799;
    ram_cell[     168] = 32'h0;  // 32'h4328a572;
    ram_cell[     169] = 32'h0;  // 32'h41dc45f4;
    ram_cell[     170] = 32'h0;  // 32'ha552c465;
    ram_cell[     171] = 32'h0;  // 32'hf1205bd9;
    ram_cell[     172] = 32'h0;  // 32'hc222bfbc;
    ram_cell[     173] = 32'h0;  // 32'h6c11e832;
    ram_cell[     174] = 32'h0;  // 32'hcb21574e;
    ram_cell[     175] = 32'h0;  // 32'h3d86def3;
    ram_cell[     176] = 32'h0;  // 32'h5a98bfe3;
    ram_cell[     177] = 32'h0;  // 32'h6baf3fc8;
    ram_cell[     178] = 32'h0;  // 32'hf3656e84;
    ram_cell[     179] = 32'h0;  // 32'h2cd7d744;
    ram_cell[     180] = 32'h0;  // 32'hb76f0e7c;
    ram_cell[     181] = 32'h0;  // 32'h8f36c7ca;
    ram_cell[     182] = 32'h0;  // 32'hca340f1f;
    ram_cell[     183] = 32'h0;  // 32'h9d5c0acc;
    ram_cell[     184] = 32'h0;  // 32'h6484c573;
    ram_cell[     185] = 32'h0;  // 32'hdeac0bc5;
    ram_cell[     186] = 32'h0;  // 32'h4f0f95bb;
    ram_cell[     187] = 32'h0;  // 32'hb20a708c;
    ram_cell[     188] = 32'h0;  // 32'hf68ae85b;
    ram_cell[     189] = 32'h0;  // 32'h0a1e2fb8;
    ram_cell[     190] = 32'h0;  // 32'ha16bc640;
    ram_cell[     191] = 32'h0;  // 32'h1ddd67df;
    ram_cell[     192] = 32'h0;  // 32'h9e28c5cb;
    ram_cell[     193] = 32'h0;  // 32'h8563fffa;
    ram_cell[     194] = 32'h0;  // 32'he7425bad;
    ram_cell[     195] = 32'h0;  // 32'h9010cd51;
    ram_cell[     196] = 32'h0;  // 32'hc3111738;
    ram_cell[     197] = 32'h0;  // 32'h56c28e07;
    ram_cell[     198] = 32'h0;  // 32'hda2ad317;
    ram_cell[     199] = 32'h0;  // 32'hfcdcbc3d;
    ram_cell[     200] = 32'h0;  // 32'hae41fc57;
    ram_cell[     201] = 32'h0;  // 32'hb8b3df7a;
    ram_cell[     202] = 32'h0;  // 32'h27006b03;
    ram_cell[     203] = 32'h0;  // 32'h6558f0ba;
    ram_cell[     204] = 32'h0;  // 32'h6e76dcbd;
    ram_cell[     205] = 32'h0;  // 32'hf4006111;
    ram_cell[     206] = 32'h0;  // 32'hadc7a1ee;
    ram_cell[     207] = 32'h0;  // 32'h050e7bbc;
    ram_cell[     208] = 32'h0;  // 32'h291518f9;
    ram_cell[     209] = 32'h0;  // 32'h26fda3f0;
    ram_cell[     210] = 32'h0;  // 32'h3cd7208b;
    ram_cell[     211] = 32'h0;  // 32'hcd39ac2e;
    ram_cell[     212] = 32'h0;  // 32'h4f57b89b;
    ram_cell[     213] = 32'h0;  // 32'hb5b2298a;
    ram_cell[     214] = 32'h0;  // 32'h63a1696e;
    ram_cell[     215] = 32'h0;  // 32'h12e8ba18;
    ram_cell[     216] = 32'h0;  // 32'h32ed079e;
    ram_cell[     217] = 32'h0;  // 32'hf0c4a725;
    ram_cell[     218] = 32'h0;  // 32'h42c72248;
    ram_cell[     219] = 32'h0;  // 32'h25a6fc32;
    ram_cell[     220] = 32'h0;  // 32'hf1d8ddb0;
    ram_cell[     221] = 32'h0;  // 32'hd9051ed9;
    ram_cell[     222] = 32'h0;  // 32'h5157c606;
    ram_cell[     223] = 32'h0;  // 32'h7924b133;
    ram_cell[     224] = 32'h0;  // 32'h66d22bdf;
    ram_cell[     225] = 32'h0;  // 32'h9de5d249;
    ram_cell[     226] = 32'h0;  // 32'h5525a33e;
    ram_cell[     227] = 32'h0;  // 32'hd8a49b92;
    ram_cell[     228] = 32'h0;  // 32'hc6ddf418;
    ram_cell[     229] = 32'h0;  // 32'hd591a183;
    ram_cell[     230] = 32'h0;  // 32'h18d66d7d;
    ram_cell[     231] = 32'h0;  // 32'h9017cbf6;
    ram_cell[     232] = 32'h0;  // 32'hfcd10507;
    ram_cell[     233] = 32'h0;  // 32'ha61a2cd7;
    ram_cell[     234] = 32'h0;  // 32'h595c60cd;
    ram_cell[     235] = 32'h0;  // 32'h0714563e;
    ram_cell[     236] = 32'h0;  // 32'hf52bd7e3;
    ram_cell[     237] = 32'h0;  // 32'hede894cd;
    ram_cell[     238] = 32'h0;  // 32'hb5dc20ed;
    ram_cell[     239] = 32'h0;  // 32'h7f222ec9;
    ram_cell[     240] = 32'h0;  // 32'h5898f495;
    ram_cell[     241] = 32'h0;  // 32'ha35228fb;
    ram_cell[     242] = 32'h0;  // 32'h7868e8cc;
    ram_cell[     243] = 32'h0;  // 32'h1d61c3de;
    ram_cell[     244] = 32'h0;  // 32'h4803dda1;
    ram_cell[     245] = 32'h0;  // 32'h913e9c44;
    ram_cell[     246] = 32'h0;  // 32'h701a1882;
    ram_cell[     247] = 32'h0;  // 32'hb2101da1;
    ram_cell[     248] = 32'h0;  // 32'hf7ee86c3;
    ram_cell[     249] = 32'h0;  // 32'h2deb9213;
    ram_cell[     250] = 32'h0;  // 32'h009f6373;
    ram_cell[     251] = 32'h0;  // 32'haff40990;
    ram_cell[     252] = 32'h0;  // 32'h092a1f03;
    ram_cell[     253] = 32'h0;  // 32'h2dc52f7c;
    ram_cell[     254] = 32'h0;  // 32'h1c6b0464;
    ram_cell[     255] = 32'h0;  // 32'hb0507aea;
    // src matrix A
    ram_cell[     256] = 32'hbd92b6b0;
    ram_cell[     257] = 32'h3bf18491;
    ram_cell[     258] = 32'h232a8adc;
    ram_cell[     259] = 32'he8a6ff97;
    ram_cell[     260] = 32'h10d1b65f;
    ram_cell[     261] = 32'h10ee65e6;
    ram_cell[     262] = 32'hfa319d71;
    ram_cell[     263] = 32'h6f45df42;
    ram_cell[     264] = 32'h39273fb1;
    ram_cell[     265] = 32'hbb501667;
    ram_cell[     266] = 32'h2ce4a709;
    ram_cell[     267] = 32'h699a7366;
    ram_cell[     268] = 32'h2e0b94e8;
    ram_cell[     269] = 32'ha3932bdb;
    ram_cell[     270] = 32'h8484878b;
    ram_cell[     271] = 32'h8feaddf3;
    ram_cell[     272] = 32'hc728756f;
    ram_cell[     273] = 32'h105be4fb;
    ram_cell[     274] = 32'hdeb8113f;
    ram_cell[     275] = 32'h7d366c79;
    ram_cell[     276] = 32'h558589f3;
    ram_cell[     277] = 32'h7ed0117d;
    ram_cell[     278] = 32'h9274504a;
    ram_cell[     279] = 32'hce30996d;
    ram_cell[     280] = 32'h7ec06aba;
    ram_cell[     281] = 32'h20e61655;
    ram_cell[     282] = 32'h902f9d45;
    ram_cell[     283] = 32'hb6f3ee7a;
    ram_cell[     284] = 32'h99c9d552;
    ram_cell[     285] = 32'h040158e3;
    ram_cell[     286] = 32'ha2334a25;
    ram_cell[     287] = 32'h62336ae9;
    ram_cell[     288] = 32'hb4e9ab12;
    ram_cell[     289] = 32'h8448a48d;
    ram_cell[     290] = 32'h2a473fd5;
    ram_cell[     291] = 32'hc37bcc5c;
    ram_cell[     292] = 32'hc094562f;
    ram_cell[     293] = 32'h8b309e2b;
    ram_cell[     294] = 32'h56f88e7e;
    ram_cell[     295] = 32'ha1bf1670;
    ram_cell[     296] = 32'hd4d029f9;
    ram_cell[     297] = 32'h00199dcd;
    ram_cell[     298] = 32'hacdcdcd6;
    ram_cell[     299] = 32'h1231e223;
    ram_cell[     300] = 32'habe4e3f4;
    ram_cell[     301] = 32'he61533c7;
    ram_cell[     302] = 32'hc008b145;
    ram_cell[     303] = 32'h7b33dad4;
    ram_cell[     304] = 32'hd1215003;
    ram_cell[     305] = 32'hcb824171;
    ram_cell[     306] = 32'hd9fdd5eb;
    ram_cell[     307] = 32'hd37bfbba;
    ram_cell[     308] = 32'h93242b5f;
    ram_cell[     309] = 32'h4a6ab8c9;
    ram_cell[     310] = 32'hfc013171;
    ram_cell[     311] = 32'hffc4f04f;
    ram_cell[     312] = 32'h502d404e;
    ram_cell[     313] = 32'h8907c58a;
    ram_cell[     314] = 32'h23a5aa03;
    ram_cell[     315] = 32'h91658d25;
    ram_cell[     316] = 32'h64d3a7ea;
    ram_cell[     317] = 32'hcac87b03;
    ram_cell[     318] = 32'h2741d5a4;
    ram_cell[     319] = 32'h8f900789;
    ram_cell[     320] = 32'h9d044cbb;
    ram_cell[     321] = 32'h48cdf6a4;
    ram_cell[     322] = 32'h148e545a;
    ram_cell[     323] = 32'h76d3f179;
    ram_cell[     324] = 32'h7fb5aedb;
    ram_cell[     325] = 32'h19538f59;
    ram_cell[     326] = 32'hc397bdd6;
    ram_cell[     327] = 32'h5de8344f;
    ram_cell[     328] = 32'h1a1afb65;
    ram_cell[     329] = 32'hed543d9a;
    ram_cell[     330] = 32'h68737b22;
    ram_cell[     331] = 32'h19a98c2c;
    ram_cell[     332] = 32'hf4513284;
    ram_cell[     333] = 32'h694ee7a5;
    ram_cell[     334] = 32'h38c3b1a1;
    ram_cell[     335] = 32'h599488dd;
    ram_cell[     336] = 32'h1d19f677;
    ram_cell[     337] = 32'ha54dbf10;
    ram_cell[     338] = 32'h3307782c;
    ram_cell[     339] = 32'h6771abb5;
    ram_cell[     340] = 32'h0feccfe8;
    ram_cell[     341] = 32'h1046674b;
    ram_cell[     342] = 32'he6b5490d;
    ram_cell[     343] = 32'h29b92337;
    ram_cell[     344] = 32'h3b3d6f43;
    ram_cell[     345] = 32'he2286f26;
    ram_cell[     346] = 32'h4a7bb918;
    ram_cell[     347] = 32'h68af2130;
    ram_cell[     348] = 32'ha6d8505f;
    ram_cell[     349] = 32'h9de502b0;
    ram_cell[     350] = 32'h96bff523;
    ram_cell[     351] = 32'hfe485c76;
    ram_cell[     352] = 32'h8a0c4b6e;
    ram_cell[     353] = 32'hb9c83bf4;
    ram_cell[     354] = 32'he2698f5e;
    ram_cell[     355] = 32'h01b30602;
    ram_cell[     356] = 32'h306aa7e4;
    ram_cell[     357] = 32'h6bec73ec;
    ram_cell[     358] = 32'hccc93204;
    ram_cell[     359] = 32'h22127a35;
    ram_cell[     360] = 32'h7ea86412;
    ram_cell[     361] = 32'hadf21471;
    ram_cell[     362] = 32'h5e101ce5;
    ram_cell[     363] = 32'h3e774447;
    ram_cell[     364] = 32'h8aea4e3d;
    ram_cell[     365] = 32'hc198ef0d;
    ram_cell[     366] = 32'h8fc23b7e;
    ram_cell[     367] = 32'hcd354ec8;
    ram_cell[     368] = 32'h1e772aa7;
    ram_cell[     369] = 32'h9d2dd805;
    ram_cell[     370] = 32'hb876359b;
    ram_cell[     371] = 32'h757c4285;
    ram_cell[     372] = 32'he0c6e215;
    ram_cell[     373] = 32'h28bbff64;
    ram_cell[     374] = 32'ha1075e7f;
    ram_cell[     375] = 32'h729f8e68;
    ram_cell[     376] = 32'hb637a876;
    ram_cell[     377] = 32'h16fe1ad4;
    ram_cell[     378] = 32'hd910f685;
    ram_cell[     379] = 32'hbb1f8c99;
    ram_cell[     380] = 32'h9fbdd086;
    ram_cell[     381] = 32'hb19dcbdb;
    ram_cell[     382] = 32'hce80e03a;
    ram_cell[     383] = 32'h3ade445e;
    ram_cell[     384] = 32'h3d27e040;
    ram_cell[     385] = 32'hc558ac37;
    ram_cell[     386] = 32'h048eaf24;
    ram_cell[     387] = 32'h2e69d254;
    ram_cell[     388] = 32'hcd7edb21;
    ram_cell[     389] = 32'h08c7bd2a;
    ram_cell[     390] = 32'h7a31c266;
    ram_cell[     391] = 32'hb8c2df29;
    ram_cell[     392] = 32'hef8833ed;
    ram_cell[     393] = 32'h493248d7;
    ram_cell[     394] = 32'hc371b348;
    ram_cell[     395] = 32'hace86503;
    ram_cell[     396] = 32'hc2a3ea33;
    ram_cell[     397] = 32'hf877876e;
    ram_cell[     398] = 32'he577d900;
    ram_cell[     399] = 32'h4f7ee719;
    ram_cell[     400] = 32'h2530362e;
    ram_cell[     401] = 32'h15e4ccbf;
    ram_cell[     402] = 32'h904ed221;
    ram_cell[     403] = 32'hbfa38eab;
    ram_cell[     404] = 32'h61e5353c;
    ram_cell[     405] = 32'h44c33d38;
    ram_cell[     406] = 32'h538f2e37;
    ram_cell[     407] = 32'h546b4f40;
    ram_cell[     408] = 32'hc7c59358;
    ram_cell[     409] = 32'h0e498bdf;
    ram_cell[     410] = 32'hcfcabd54;
    ram_cell[     411] = 32'h9dd05cc2;
    ram_cell[     412] = 32'h303e7a1c;
    ram_cell[     413] = 32'ha3849565;
    ram_cell[     414] = 32'hd93c2c7e;
    ram_cell[     415] = 32'h721a748a;
    ram_cell[     416] = 32'h3a4b8d4c;
    ram_cell[     417] = 32'hfa561a13;
    ram_cell[     418] = 32'h04edefbb;
    ram_cell[     419] = 32'h2770cf20;
    ram_cell[     420] = 32'h9347fe4f;
    ram_cell[     421] = 32'ha7307771;
    ram_cell[     422] = 32'hbd7e6b68;
    ram_cell[     423] = 32'h0839d094;
    ram_cell[     424] = 32'h86de6922;
    ram_cell[     425] = 32'h237449dc;
    ram_cell[     426] = 32'hebff999c;
    ram_cell[     427] = 32'h1010faa9;
    ram_cell[     428] = 32'he70aa227;
    ram_cell[     429] = 32'h5d3e704f;
    ram_cell[     430] = 32'hd412a079;
    ram_cell[     431] = 32'h42122f30;
    ram_cell[     432] = 32'hcef25c7d;
    ram_cell[     433] = 32'hb3043a96;
    ram_cell[     434] = 32'h7a02a158;
    ram_cell[     435] = 32'hd46b1d88;
    ram_cell[     436] = 32'hd4160db4;
    ram_cell[     437] = 32'h538afab0;
    ram_cell[     438] = 32'h140fb509;
    ram_cell[     439] = 32'h4d99eafd;
    ram_cell[     440] = 32'h77925ecc;
    ram_cell[     441] = 32'h6436ff4d;
    ram_cell[     442] = 32'h209e105f;
    ram_cell[     443] = 32'h95bd6540;
    ram_cell[     444] = 32'h44b42fa4;
    ram_cell[     445] = 32'h07358559;
    ram_cell[     446] = 32'h3bbaab44;
    ram_cell[     447] = 32'hbba08383;
    ram_cell[     448] = 32'h935a3627;
    ram_cell[     449] = 32'h37da93e0;
    ram_cell[     450] = 32'h444d4859;
    ram_cell[     451] = 32'h84487e74;
    ram_cell[     452] = 32'h0aeeca07;
    ram_cell[     453] = 32'h15d547cc;
    ram_cell[     454] = 32'hcc7cf01a;
    ram_cell[     455] = 32'h95ae153f;
    ram_cell[     456] = 32'ha6352e4c;
    ram_cell[     457] = 32'hd74c72f0;
    ram_cell[     458] = 32'hd514d138;
    ram_cell[     459] = 32'he616667f;
    ram_cell[     460] = 32'hf0ce410f;
    ram_cell[     461] = 32'hb5f2da03;
    ram_cell[     462] = 32'h1aeb5ac6;
    ram_cell[     463] = 32'h235f1bd5;
    ram_cell[     464] = 32'hec7038d3;
    ram_cell[     465] = 32'hcde54275;
    ram_cell[     466] = 32'hedf784e3;
    ram_cell[     467] = 32'hdea34200;
    ram_cell[     468] = 32'h47c63197;
    ram_cell[     469] = 32'hade06ae0;
    ram_cell[     470] = 32'hdf254081;
    ram_cell[     471] = 32'hb1f1be8b;
    ram_cell[     472] = 32'hd8d38e43;
    ram_cell[     473] = 32'h5e447afd;
    ram_cell[     474] = 32'h6075cff6;
    ram_cell[     475] = 32'h99d0ba92;
    ram_cell[     476] = 32'h0da7ad8d;
    ram_cell[     477] = 32'h562da6ca;
    ram_cell[     478] = 32'he28f742d;
    ram_cell[     479] = 32'h1bfa367e;
    ram_cell[     480] = 32'h77c79028;
    ram_cell[     481] = 32'h75d3ed7b;
    ram_cell[     482] = 32'h39492851;
    ram_cell[     483] = 32'hf470160b;
    ram_cell[     484] = 32'hbb141ee6;
    ram_cell[     485] = 32'hadbbb97b;
    ram_cell[     486] = 32'ha3543a49;
    ram_cell[     487] = 32'h4af123e7;
    ram_cell[     488] = 32'hd37027bb;
    ram_cell[     489] = 32'h6da29309;
    ram_cell[     490] = 32'h7d8a73de;
    ram_cell[     491] = 32'hdca2a5d1;
    ram_cell[     492] = 32'h1115c7b0;
    ram_cell[     493] = 32'h6044fb36;
    ram_cell[     494] = 32'h32e09e8f;
    ram_cell[     495] = 32'h53baeea2;
    ram_cell[     496] = 32'h946976de;
    ram_cell[     497] = 32'h1d93ca06;
    ram_cell[     498] = 32'h35f1df44;
    ram_cell[     499] = 32'h37093464;
    ram_cell[     500] = 32'h6315c22d;
    ram_cell[     501] = 32'h711c2d83;
    ram_cell[     502] = 32'h101f2f6c;
    ram_cell[     503] = 32'he7e8afbc;
    ram_cell[     504] = 32'h6ae4ce98;
    ram_cell[     505] = 32'h560d1ba5;
    ram_cell[     506] = 32'h53dffc7a;
    ram_cell[     507] = 32'h12ded174;
    ram_cell[     508] = 32'h17073a2e;
    ram_cell[     509] = 32'hf2d87998;
    ram_cell[     510] = 32'hb02e228d;
    ram_cell[     511] = 32'h273ca35b;
    // src matrix B
    ram_cell[     512] = 32'hdb871783;
    ram_cell[     513] = 32'ha1975928;
    ram_cell[     514] = 32'hf26f0983;
    ram_cell[     515] = 32'h91f78334;
    ram_cell[     516] = 32'h9c967bec;
    ram_cell[     517] = 32'hd3844973;
    ram_cell[     518] = 32'h044645c9;
    ram_cell[     519] = 32'h118157d4;
    ram_cell[     520] = 32'h6f912af5;
    ram_cell[     521] = 32'hdf8236a9;
    ram_cell[     522] = 32'h8954dab9;
    ram_cell[     523] = 32'h5e9b23a9;
    ram_cell[     524] = 32'h1051097d;
    ram_cell[     525] = 32'h62c70a70;
    ram_cell[     526] = 32'h66eb2254;
    ram_cell[     527] = 32'hb2f0560e;
    ram_cell[     528] = 32'h7432d563;
    ram_cell[     529] = 32'h464e8620;
    ram_cell[     530] = 32'h8fc2453c;
    ram_cell[     531] = 32'he0611ed8;
    ram_cell[     532] = 32'h5cf6a717;
    ram_cell[     533] = 32'h49b675c9;
    ram_cell[     534] = 32'h3002185f;
    ram_cell[     535] = 32'h72fd4f71;
    ram_cell[     536] = 32'hc931e381;
    ram_cell[     537] = 32'habd6c842;
    ram_cell[     538] = 32'hfde4ad1a;
    ram_cell[     539] = 32'he4e60527;
    ram_cell[     540] = 32'ha0b67fa0;
    ram_cell[     541] = 32'h1f6c537e;
    ram_cell[     542] = 32'h1443a682;
    ram_cell[     543] = 32'h7eef1e19;
    ram_cell[     544] = 32'he8d3862c;
    ram_cell[     545] = 32'h8c454860;
    ram_cell[     546] = 32'h9c525373;
    ram_cell[     547] = 32'hb2b5dc44;
    ram_cell[     548] = 32'ha531177a;
    ram_cell[     549] = 32'hc718947a;
    ram_cell[     550] = 32'h6195fe69;
    ram_cell[     551] = 32'ha5e6cbb5;
    ram_cell[     552] = 32'h88e26e4f;
    ram_cell[     553] = 32'hb642aa38;
    ram_cell[     554] = 32'hdf234235;
    ram_cell[     555] = 32'h34c84b35;
    ram_cell[     556] = 32'h46df617d;
    ram_cell[     557] = 32'h7ae6bef0;
    ram_cell[     558] = 32'hc5b14ce5;
    ram_cell[     559] = 32'ha8f2a4b5;
    ram_cell[     560] = 32'he3c3e5ef;
    ram_cell[     561] = 32'h2807550c;
    ram_cell[     562] = 32'h94a6227d;
    ram_cell[     563] = 32'hb5075982;
    ram_cell[     564] = 32'h124af2c3;
    ram_cell[     565] = 32'h7a6fa558;
    ram_cell[     566] = 32'h8ca88e03;
    ram_cell[     567] = 32'ha305f294;
    ram_cell[     568] = 32'h18ed919d;
    ram_cell[     569] = 32'he089aeab;
    ram_cell[     570] = 32'hd0462d2a;
    ram_cell[     571] = 32'hd5e04713;
    ram_cell[     572] = 32'hb3ad6ce0;
    ram_cell[     573] = 32'h61c90eb0;
    ram_cell[     574] = 32'h981f38fd;
    ram_cell[     575] = 32'he9fc8a4c;
    ram_cell[     576] = 32'h199e7c07;
    ram_cell[     577] = 32'hed34b5a4;
    ram_cell[     578] = 32'hbe682490;
    ram_cell[     579] = 32'h2e056969;
    ram_cell[     580] = 32'h599fdddc;
    ram_cell[     581] = 32'h26ead1a4;
    ram_cell[     582] = 32'h74cb7680;
    ram_cell[     583] = 32'h1eebd482;
    ram_cell[     584] = 32'h18dd3d0f;
    ram_cell[     585] = 32'h9f436e41;
    ram_cell[     586] = 32'h2b08ede8;
    ram_cell[     587] = 32'h2c43a8eb;
    ram_cell[     588] = 32'h3b18f33e;
    ram_cell[     589] = 32'h3a42ae78;
    ram_cell[     590] = 32'h7d32f1e6;
    ram_cell[     591] = 32'hc4840d55;
    ram_cell[     592] = 32'h3a4f9d26;
    ram_cell[     593] = 32'he4257d66;
    ram_cell[     594] = 32'hfe364a8a;
    ram_cell[     595] = 32'h0dc0c49e;
    ram_cell[     596] = 32'h73622f5e;
    ram_cell[     597] = 32'h5bd7dc78;
    ram_cell[     598] = 32'hfa2bfda6;
    ram_cell[     599] = 32'h50467d8f;
    ram_cell[     600] = 32'hb12edf92;
    ram_cell[     601] = 32'hf64612b2;
    ram_cell[     602] = 32'h31d10fd6;
    ram_cell[     603] = 32'hc2794186;
    ram_cell[     604] = 32'h8ac1945e;
    ram_cell[     605] = 32'h6baf04d4;
    ram_cell[     606] = 32'hefaf4806;
    ram_cell[     607] = 32'h4dece29c;
    ram_cell[     608] = 32'hc2342875;
    ram_cell[     609] = 32'h9024a4bf;
    ram_cell[     610] = 32'hd01982e2;
    ram_cell[     611] = 32'h252d2683;
    ram_cell[     612] = 32'had3360b6;
    ram_cell[     613] = 32'h05b031f4;
    ram_cell[     614] = 32'h67ed3e93;
    ram_cell[     615] = 32'hfdad8812;
    ram_cell[     616] = 32'h23b64c17;
    ram_cell[     617] = 32'he2c6eb51;
    ram_cell[     618] = 32'h8aea9c28;
    ram_cell[     619] = 32'h8c717e94;
    ram_cell[     620] = 32'hb1213d9d;
    ram_cell[     621] = 32'h475dcbd2;
    ram_cell[     622] = 32'h4ff44f34;
    ram_cell[     623] = 32'h4edac10b;
    ram_cell[     624] = 32'hc4b0abe7;
    ram_cell[     625] = 32'hb5333664;
    ram_cell[     626] = 32'h1d9c722e;
    ram_cell[     627] = 32'hc10870ff;
    ram_cell[     628] = 32'h6c6e924e;
    ram_cell[     629] = 32'h3a70ebc9;
    ram_cell[     630] = 32'h8fc69a29;
    ram_cell[     631] = 32'h8af62e40;
    ram_cell[     632] = 32'h0906115d;
    ram_cell[     633] = 32'h9430b792;
    ram_cell[     634] = 32'hdb3914fd;
    ram_cell[     635] = 32'hdad65a4f;
    ram_cell[     636] = 32'h93564246;
    ram_cell[     637] = 32'h850a957f;
    ram_cell[     638] = 32'h8b648d35;
    ram_cell[     639] = 32'hda929163;
    ram_cell[     640] = 32'h3ae97512;
    ram_cell[     641] = 32'h422b143a;
    ram_cell[     642] = 32'h1fd2e1d0;
    ram_cell[     643] = 32'h8d359478;
    ram_cell[     644] = 32'hfab75d36;
    ram_cell[     645] = 32'hf8bca1db;
    ram_cell[     646] = 32'h78c99464;
    ram_cell[     647] = 32'h61c33fbd;
    ram_cell[     648] = 32'h4c8326da;
    ram_cell[     649] = 32'h83772afd;
    ram_cell[     650] = 32'hb7a6eb3f;
    ram_cell[     651] = 32'hca35e4c7;
    ram_cell[     652] = 32'h245d94e8;
    ram_cell[     653] = 32'hd6021b33;
    ram_cell[     654] = 32'hc636e70f;
    ram_cell[     655] = 32'hdc756fae;
    ram_cell[     656] = 32'h268dc6e7;
    ram_cell[     657] = 32'h03d68ce3;
    ram_cell[     658] = 32'h853d93ae;
    ram_cell[     659] = 32'ha84196ce;
    ram_cell[     660] = 32'h29a6227d;
    ram_cell[     661] = 32'ha0b1b763;
    ram_cell[     662] = 32'h4f77f5fd;
    ram_cell[     663] = 32'hbc71cef4;
    ram_cell[     664] = 32'h75d7fc34;
    ram_cell[     665] = 32'h5f932b4d;
    ram_cell[     666] = 32'he575ff07;
    ram_cell[     667] = 32'h250d3a21;
    ram_cell[     668] = 32'h60612d73;
    ram_cell[     669] = 32'h8c228016;
    ram_cell[     670] = 32'h06c1a715;
    ram_cell[     671] = 32'hfe56aa6c;
    ram_cell[     672] = 32'hbc6cb460;
    ram_cell[     673] = 32'hee607d9f;
    ram_cell[     674] = 32'h9ba95d4d;
    ram_cell[     675] = 32'h7e6a4604;
    ram_cell[     676] = 32'h4d30be77;
    ram_cell[     677] = 32'h9df44176;
    ram_cell[     678] = 32'h45f97a88;
    ram_cell[     679] = 32'h9855d307;
    ram_cell[     680] = 32'h8d36e51b;
    ram_cell[     681] = 32'h97ee627d;
    ram_cell[     682] = 32'h548a669e;
    ram_cell[     683] = 32'haa3976a4;
    ram_cell[     684] = 32'hf08f0cdf;
    ram_cell[     685] = 32'h3543dd05;
    ram_cell[     686] = 32'hcaad9034;
    ram_cell[     687] = 32'hdb39d761;
    ram_cell[     688] = 32'had7e4435;
    ram_cell[     689] = 32'h3cdc498e;
    ram_cell[     690] = 32'hcd194b0c;
    ram_cell[     691] = 32'h409396f8;
    ram_cell[     692] = 32'h78c35209;
    ram_cell[     693] = 32'hfbd8e722;
    ram_cell[     694] = 32'h11b387c8;
    ram_cell[     695] = 32'hae1d7ebe;
    ram_cell[     696] = 32'h60cebdc6;
    ram_cell[     697] = 32'hc1d112ee;
    ram_cell[     698] = 32'h332f6965;
    ram_cell[     699] = 32'h80ca7413;
    ram_cell[     700] = 32'h9821ba64;
    ram_cell[     701] = 32'hd2cd2091;
    ram_cell[     702] = 32'h315c147a;
    ram_cell[     703] = 32'haf67a444;
    ram_cell[     704] = 32'h1dd4cfd0;
    ram_cell[     705] = 32'hbc68cd3f;
    ram_cell[     706] = 32'h040e072f;
    ram_cell[     707] = 32'he0a940e7;
    ram_cell[     708] = 32'h076eaf85;
    ram_cell[     709] = 32'hdf979526;
    ram_cell[     710] = 32'h2fc03181;
    ram_cell[     711] = 32'h1ca109ad;
    ram_cell[     712] = 32'hfb002616;
    ram_cell[     713] = 32'hac21411b;
    ram_cell[     714] = 32'hde6f8da9;
    ram_cell[     715] = 32'hdcca6002;
    ram_cell[     716] = 32'h08a95096;
    ram_cell[     717] = 32'hd44a4903;
    ram_cell[     718] = 32'hdc526ac4;
    ram_cell[     719] = 32'h5bf0ff1f;
    ram_cell[     720] = 32'h650bee03;
    ram_cell[     721] = 32'h168434f8;
    ram_cell[     722] = 32'hbcee1678;
    ram_cell[     723] = 32'h10f3b3b5;
    ram_cell[     724] = 32'h42fe6f06;
    ram_cell[     725] = 32'hb69ee61b;
    ram_cell[     726] = 32'h3905e353;
    ram_cell[     727] = 32'haf479fdb;
    ram_cell[     728] = 32'h3d6ad593;
    ram_cell[     729] = 32'h30c388a5;
    ram_cell[     730] = 32'hbb287052;
    ram_cell[     731] = 32'h04b39d54;
    ram_cell[     732] = 32'hae39bd8b;
    ram_cell[     733] = 32'h031c469e;
    ram_cell[     734] = 32'hef93cd5f;
    ram_cell[     735] = 32'heeeb6a02;
    ram_cell[     736] = 32'he799225b;
    ram_cell[     737] = 32'ha7d3d9fb;
    ram_cell[     738] = 32'h5dafc0c6;
    ram_cell[     739] = 32'hbd6f320e;
    ram_cell[     740] = 32'h22edf72c;
    ram_cell[     741] = 32'hb81bebf1;
    ram_cell[     742] = 32'hafac0c9f;
    ram_cell[     743] = 32'h4e4c1466;
    ram_cell[     744] = 32'hed88ac18;
    ram_cell[     745] = 32'ha85b6819;
    ram_cell[     746] = 32'hd725f554;
    ram_cell[     747] = 32'he3920a75;
    ram_cell[     748] = 32'ha1f987c2;
    ram_cell[     749] = 32'h3507d3ae;
    ram_cell[     750] = 32'h5385d61c;
    ram_cell[     751] = 32'h95c4c2d3;
    ram_cell[     752] = 32'hac73c368;
    ram_cell[     753] = 32'h67cc1c13;
    ram_cell[     754] = 32'h3b0d8b4e;
    ram_cell[     755] = 32'h7fb3d9d1;
    ram_cell[     756] = 32'h2b60125e;
    ram_cell[     757] = 32'h7453be5c;
    ram_cell[     758] = 32'h064badc0;
    ram_cell[     759] = 32'h6ee90bac;
    ram_cell[     760] = 32'h3ec30de0;
    ram_cell[     761] = 32'hdbd4710a;
    ram_cell[     762] = 32'hcd453dd0;
    ram_cell[     763] = 32'hbd974cdf;
    ram_cell[     764] = 32'h075443f0;
    ram_cell[     765] = 32'h5ef90078;
    ram_cell[     766] = 32'h1f8ee097;
    ram_cell[     767] = 32'hdcf6fe08;
end

endmodule
